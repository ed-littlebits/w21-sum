CircuitMaker Text
5.6
Probes: 5
U2D_14
AC Analysis
0 504 415 65280
U2D_14
Transient Analysis
0 505 423 65280
U2D_1
Operating Point
0 503 449 65280
vs1#branch
DC Sweep
0 167 289 65280
U2D_1
Transfer Function
0 505 448 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
10 180 30 240 10
1542 -237 3284 747
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 2 0
20 Package,Description,
48 C:\Program Files\CircuitMaker 2000 Trial\BOM.DAT
5 7
3 4 0.328025 0.500000
1542 -237 2413 747
77070354 336
2
2 

2 

0
0
0
32
9 V Source~
197 184 288 0 2 5
0 13 6
0
0 0 17264 90
1 0
-4 -20 3 -12
3 Vs1
-8 -30 13 -22
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
9429 0 0
2
41646.5 0
0
11 Signal Gen~
195 41 208 0 64 64
0 9 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 1075838976 1065353216
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 264
20
1 1000 2.5 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
8 1.5/3.5V
-28 -30 28 -22
2 V2
-7 -40 7 -32
0
0
38 %D %1 %2 DC 0 SIN(2.5 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
7437 0 0
2
41646.4 0
0
11 Signal Gen~
195 39 383 0 19 64
0 8 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1149861888 1075838976 1065353216
20
1 1100 2.5 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
8 1.5/3.5V
-29 -30 27 -22
2 V1
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 SIN(2.5 1 1.1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
6197 0 0
2
41646.4 0
0
7 Ground~
168 440 359 0 1 3
0 2
0
0 0 53360 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7170 0 0
2
41646.4 1
0
10 Capacitor~
219 440 330 0 2 5
0 2 3
0
0 0 848 90
3 .1u
11 0 32 8
2 C4
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3938 0 0
2
41646.4 0
0
7 Ground~
168 376 417 0 1 3
0 2
0
0 0 53360 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7781 0 0
2
41646.4 0
0
9 Terminal~
194 456 419 0 1 3
0 3
0
0 0 49520 0
4 vpos
-14 -13 14 -5
2 T5
-7 -32 7 -24
0
5 vpos;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5978 0 0
2
41646.4 2
0
7 Ground~
168 456 476 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9486 0 0
2
41646.4 1
0
8 Op-Amp5~
219 456 450 0 5 11
0 11 7 3 2 10
0
0 0 848 0
10 LM6132A/NS
16 11 86 19
3 U2D
18 23 39 31
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
5 SMD8A
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 62
88 0 0 256 2 1 3 0
1 U
5847 0 0
2
41646.4 0
0
7 Ground~
168 166 535 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3503 0 0
2
41646.4 8
0
8 Op-Amp5~
219 222 457 0 5 11
0 12 4 3 2 4
0
0 0 848 0
10 LM6132A/NS
14 24 84 32
3 U1B
27 8 48 16
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
5 SMD8A
16

0 5 6 8 4 7 3 2 8 4
1 5 6 8 4 7 50
88 0 0 256 2 2 2 0
1 U
3983 0 0
2
41646.4 7
0
7 Ground~
168 222 477 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
858 0 0
2
41646.4 6
0
9 Terminal~
194 222 427 0 1 3
0 3
0
0 0 49520 0
4 vpos
-14 -13 14 -5
2 T4
-7 -32 7 -24
0
5 vpos;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6251 0 0
2
41646.4 5
0
10 Capacitor~
219 82 465 0 2 5
0 2 3
0
0 0 848 90
3 .1u
11 0 32 8
2 C3
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
384 0 0
2
41646.4 2
0
7 Ground~
168 82 494 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4542 0 0
2
41646.4 1
0
9 Terminal~
194 83 437 0 1 3
0 3
0
0 0 49520 0
4 vpos
-14 -13 14 -5
2 T2
-7 -32 7 -24
0
5 vpos;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3308 0 0
2
41646.4 0
0
9 Terminal~
194 86 256 0 1 3
0 3
0
0 0 49520 0
4 vpos
-14 -13 14 -5
2 T1
-7 -32 7 -24
0
5 vpos;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3355 0 0
2
41646.4 0
0
7 Ground~
168 86 319 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5771 0 0
2
41646.4 0
0
10 Capacitor~
219 87 288 0 2 5
0 2 3
0
0 0 848 90
3 .1u
11 0 32 8
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3200 0 0
2
41646.4 0
0
2 +V
167 440 304 0 1 3
0 3
0
0 0 54640 0
2 5V
9 -6 23 2
2 V4
-7 -32 7 -24
4 vpos
-39 -7 -11 1
5 vpos;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3494 0 0
2
5.89614e-315 0
0
9 Terminal~
194 226 252 0 1 3
0 3
0
0 0 49520 0
4 vpos
-14 -13 14 -5
2 T3
-7 -32 7 -24
0
5 vpos;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6920 0 0
2
5.89614e-315 5.46559e-315
0
7 Ground~
168 226 302 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6534 0 0
2
5.89614e-315 5.46041e-315
0
8 Op-Amp5~
219 226 282 0 5 11
0 6 5 3 2 5
0
0 0 848 0
10 LM6132A/NS
19 10 89 18
3 U1A
43 0 64 8
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
5 SMD8A
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 70
88 0 0 256 2 1 2 0
1 U
810 0 0
2
5.89614e-315 5.45782e-315
0
7 Ground~
168 170 360 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5116 0 0
2
5.89614e-315 5.34643e-315
0
9 Resistor~
219 400 399 0 3 5
0 2 7 -1
0
0 0 880 0
4 100k
-13 -14 15 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4787 0 0
2
41646.4 0
0
9 Resistor~
219 486 399 0 2 5
0 7 10
0
0 0 880 0
4 200k
-12 -14 16 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5926 0 0
2
41646.4 0
0
9 Resistor~
219 292 457 0 2 5
0 4 11
0
0 0 880 0
4 100k
-12 -14 16 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4713 0 0
2
41646.4 10
0
9 Resistor~
219 152 427 0 2 5
0 12 8
0
0 0 880 90
4 100k
-34 3 -6 11
2 R2
-24 -11 -10 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6623 0 0
2
41646.4 9
0
9 Resistor~
219 153 502 0 3 5
0 2 12 -1
0
0 0 880 90
4 200k
-34 3 -6 11
2 R1
-24 -11 -10 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3120 0 0
2
41646.4 3
0
9 Resistor~
219 157 327 0 3 5
0 2 13 -1
0
0 0 880 90
4 200k
-34 3 -6 11
3 R23
-27 -11 -6 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5649 0 0
2
41646.4 0
0
9 Resistor~
219 156 252 0 2 5
0 13 9
0
0 0 880 90
4 100k
-34 3 -6 11
2 R8
-24 -11 -10 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6227 0 0
2
5.89614e-315 5.49149e-315
0
9 Resistor~
219 296 282 0 2 5
0 5 11
0
0 0 880 0
4 100k
-12 -14 16 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3426 0 0
2
5.89614e-315 5.47207e-315
0
33
1 0 4 0 0 4096 0 27 0 0 5 2
274 457
248 457
2 0 5 0 0 8320 0 23 0 0 30 4
208 276
208 235
261 235
261 282
2 1 6 0 0 4224 0 1 23 0 0 2
205 288
208 288
2 0 7 0 0 8192 0 9 0 0 14 3
438 444
428 444
428 399
5 2 4 0 0 12416 0 11 11 0 0 6
240 457
248 457
248 406
189 406
189 451
204 451
2 1 2 0 0 16512 0 2 18 0 0 6
72 213
84 213
84 235
50 235
50 313
86 313
2 0 2 0 0 0 0 3 0 0 20 5
70 388
70 417
49 417
49 483
82 483
1 2 8 0 0 4224 0 3 28 0 0 3
70 378
152 378
152 409
1 2 9 0 0 4224 0 2 31 0 0 3
72 203
156 203
156 234
1 2 3 0 0 4096 0 20 5 0 0 2
440 313
440 321
1 1 2 0 0 0 0 4 5 0 0 2
440 353
440 339
5 2 10 0 0 8320 0 9 26 0 0 3
474 450
504 450
504 399
1 1 2 0 0 16 0 6 25 0 0 3
376 411
376 399
382 399
2 1 7 0 0 4224 0 25 26 0 0 2
418 399
468 399
2 0 11 0 0 8192 0 27 0 0 16 3
310 457
310 456
338 456
2 1 11 0 0 8320 0 32 9 0 0 4
314 282
338 282
338 456
438 456
1 3 3 0 0 4096 0 7 9 0 0 4
456 428
456 440
456 440
456 437
4 1 2 0 0 0 0 9 8 0 0 2
456 463
456 470
1 2 3 0 0 0 0 16 14 0 0 3
83 446
83 456
82 456
1 1 2 0 0 0 0 15 14 0 0 2
82 488
82 474
1 1 2 0 0 0 0 10 29 0 0 3
166 529
166 520
153 520
2 0 12 0 0 4096 0 29 0 0 23 3
153 484
153 463
152 463
1 1 12 0 0 8320 0 28 11 0 0 3
152 445
152 463
204 463
1 3 3 0 0 0 0 13 11 0 0 2
222 436
222 444
4 1 2 0 0 0 0 11 12 0 0 2
222 470
222 471
1 2 3 0 0 8320 0 17 19 0 0 3
86 265
87 265
87 279
1 1 2 0 0 0 0 18 19 0 0 4
86 313
86 306
87 306
87 297
1 1 2 0 0 0 0 24 30 0 0 3
170 354
170 345
157 345
2 0 13 0 0 4224 0 30 0 0 31 3
157 309
157 288
156 288
1 5 5 0 0 0 0 32 23 0 0 2
278 282
244 282
1 1 13 0 0 128 0 31 1 0 0 3
156 270
156 288
163 288
1 3 3 0 0 0 0 21 23 0 0 2
226 261
226 269
4 1 2 0 0 0 0 23 22 0 0 2
226 295
226 296
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
425 182 480 226
428 184 476 216
6 notes:
0
2 0 0
2 V2
0
2 V1
2 2.5 0.5
2 V2
0.5 1 0.5
100 1 1 1e+06
0 0.005 2e-05 2e-05
0
0
0 0 0
0 0 0
2 V2
0
10 0 1 20
0
0 0 0 0 0
14208 10 40 10
2 R7
0.001 51000 12500
2 r9
0.001 51000 12500
100 -1 1 20 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
